-- system.vhd

-- Generated using ACDS version 17.1 590

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;

entity system is
	port (
		audio_codec_external_interface_ADCDAT  : in    std_logic := '0'; --  audio_codec_external_interface.ADCDAT
		audio_codec_external_interface_ADCLRCK : in    std_logic := '0'; --                                .ADCLRCK
		audio_codec_external_interface_BCLK    : in    std_logic := '0'; --                                .BCLK
		audio_codec_external_interface_DACDAT  : out   std_logic;        --                                .DACDAT
		audio_codec_external_interface_DACLRCK : in    std_logic := '0'; --                                .DACLRCK
		audio_config_external_interface_SDAT   : inout std_logic := '0'; -- audio_config_external_interface.SDAT
		audio_config_external_interface_SCLK   : out   std_logic;        --                                .SCLK
		audio_pll_1_audio_clk_clk              : out   std_logic;        --           audio_pll_1_audio_clk.clk
		clk_clk                                : in    std_logic := '0'; --                             clk.clk
		reset_reset_n                          : in    std_logic := '0'  --                           reset.reset_n
	);
end entity system;

architecture rtl of system is
	component system_audio_codec is
		port (
			clk         : in  std_logic                     := 'X';             -- clk
			reset       : in  std_logic                     := 'X';             -- reset
			address     : in  std_logic_vector(1 downto 0)  := (others => 'X'); -- address
			chipselect  : in  std_logic                     := 'X';             -- chipselect
			read        : in  std_logic                     := 'X';             -- read
			write       : in  std_logic                     := 'X';             -- write
			writedata   : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			readdata    : out std_logic_vector(31 downto 0);                    -- readdata
			irq         : out std_logic;                                        -- irq
			AUD_ADCDAT  : in  std_logic                     := 'X';             -- export
			AUD_ADCLRCK : in  std_logic                     := 'X';             -- export
			AUD_BCLK    : in  std_logic                     := 'X';             -- export
			AUD_DACDAT  : out std_logic;                                        -- export
			AUD_DACLRCK : in  std_logic                     := 'X'              -- export
		);
	end component system_audio_codec;

	component system_audio_config is
		port (
			clk         : in    std_logic                     := 'X';             -- clk
			reset       : in    std_logic                     := 'X';             -- reset
			address     : in    std_logic_vector(1 downto 0)  := (others => 'X'); -- address
			byteenable  : in    std_logic_vector(3 downto 0)  := (others => 'X'); -- byteenable
			read        : in    std_logic                     := 'X';             -- read
			write       : in    std_logic                     := 'X';             -- write
			writedata   : in    std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			readdata    : out   std_logic_vector(31 downto 0);                    -- readdata
			waitrequest : out   std_logic;                                        -- waitrequest
			I2C_SDAT    : inout std_logic                     := 'X';             -- export
			I2C_SCLK    : out   std_logic                                         -- export
		);
	end component system_audio_config;

	component system_audio_pll_0 is
		port (
			ref_clk_clk        : in  std_logic := 'X'; -- clk
			ref_reset_reset    : in  std_logic := 'X'; -- reset
			audio_clk_clk      : out std_logic;        -- clk
			reset_source_reset : out std_logic         -- reset
		);
	end component system_audio_pll_0;

	component system_nios2_gen2_0 is
		port (
			clk                                 : in  std_logic                     := 'X';             -- clk
			reset_n                             : in  std_logic                     := 'X';             -- reset_n
			reset_req                           : in  std_logic                     := 'X';             -- reset_req
			d_address                           : out std_logic_vector(20 downto 0);                    -- address
			d_byteenable                        : out std_logic_vector(3 downto 0);                     -- byteenable
			d_read                              : out std_logic;                                        -- read
			d_readdata                          : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			d_waitrequest                       : in  std_logic                     := 'X';             -- waitrequest
			d_write                             : out std_logic;                                        -- write
			d_writedata                         : out std_logic_vector(31 downto 0);                    -- writedata
			debug_mem_slave_debugaccess_to_roms : out std_logic;                                        -- debugaccess
			i_address                           : out std_logic_vector(20 downto 0);                    -- address
			i_read                              : out std_logic;                                        -- read
			i_readdata                          : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			i_waitrequest                       : in  std_logic                     := 'X';             -- waitrequest
			irq                                 : in  std_logic_vector(31 downto 0) := (others => 'X'); -- irq
			debug_reset_request                 : out std_logic;                                        -- reset
			debug_mem_slave_address             : in  std_logic_vector(8 downto 0)  := (others => 'X'); -- address
			debug_mem_slave_byteenable          : in  std_logic_vector(3 downto 0)  := (others => 'X'); -- byteenable
			debug_mem_slave_debugaccess         : in  std_logic                     := 'X';             -- debugaccess
			debug_mem_slave_read                : in  std_logic                     := 'X';             -- read
			debug_mem_slave_readdata            : out std_logic_vector(31 downto 0);                    -- readdata
			debug_mem_slave_waitrequest         : out std_logic;                                        -- waitrequest
			debug_mem_slave_write               : in  std_logic                     := 'X';             -- write
			debug_mem_slave_writedata           : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			dummy_ci_port                       : out std_logic                                         -- readra
		);
	end component system_nios2_gen2_0;

	component system_onchip_memory2_0 is
		port (
			clk        : in  std_logic                     := 'X';             -- clk
			address    : in  std_logic_vector(16 downto 0) := (others => 'X'); -- address
			clken      : in  std_logic                     := 'X';             -- clken
			chipselect : in  std_logic                     := 'X';             -- chipselect
			write      : in  std_logic                     := 'X';             -- write
			readdata   : out std_logic_vector(31 downto 0);                    -- readdata
			writedata  : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			byteenable : in  std_logic_vector(3 downto 0)  := (others => 'X'); -- byteenable
			reset      : in  std_logic                     := 'X';             -- reset
			reset_req  : in  std_logic                     := 'X';             -- reset_req
			freeze     : in  std_logic                     := 'X'              -- freeze
		);
	end component system_onchip_memory2_0;

	component system_sysid_qsys_0 is
		port (
			clock    : in  std_logic                     := 'X'; -- clk
			reset_n  : in  std_logic                     := 'X'; -- reset_n
			readdata : out std_logic_vector(31 downto 0);        -- readdata
			address  : in  std_logic                     := 'X'  -- address
		);
	end component system_sysid_qsys_0;

	component system_mm_interconnect_0 is
		port (
			clk_0_clk_clk                                   : in  std_logic                     := 'X';             -- clk
			clock_bridge_0_out_clk_clk                      : in  std_logic                     := 'X';             -- clk
			audio_codec_reset_reset_bridge_in_reset_reset   : in  std_logic                     := 'X';             -- reset
			nios2_gen2_0_reset_reset_bridge_in_reset_reset  : in  std_logic                     := 'X';             -- reset
			nios2_gen2_0_data_master_address                : in  std_logic_vector(20 downto 0) := (others => 'X'); -- address
			nios2_gen2_0_data_master_waitrequest            : out std_logic;                                        -- waitrequest
			nios2_gen2_0_data_master_byteenable             : in  std_logic_vector(3 downto 0)  := (others => 'X'); -- byteenable
			nios2_gen2_0_data_master_read                   : in  std_logic                     := 'X';             -- read
			nios2_gen2_0_data_master_readdata               : out std_logic_vector(31 downto 0);                    -- readdata
			nios2_gen2_0_data_master_write                  : in  std_logic                     := 'X';             -- write
			nios2_gen2_0_data_master_writedata              : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			nios2_gen2_0_data_master_debugaccess            : in  std_logic                     := 'X';             -- debugaccess
			nios2_gen2_0_instruction_master_address         : in  std_logic_vector(20 downto 0) := (others => 'X'); -- address
			nios2_gen2_0_instruction_master_waitrequest     : out std_logic;                                        -- waitrequest
			nios2_gen2_0_instruction_master_read            : in  std_logic                     := 'X';             -- read
			nios2_gen2_0_instruction_master_readdata        : out std_logic_vector(31 downto 0);                    -- readdata
			audio_codec_avalon_audio_slave_address          : out std_logic_vector(1 downto 0);                     -- address
			audio_codec_avalon_audio_slave_write            : out std_logic;                                        -- write
			audio_codec_avalon_audio_slave_read             : out std_logic;                                        -- read
			audio_codec_avalon_audio_slave_readdata         : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			audio_codec_avalon_audio_slave_writedata        : out std_logic_vector(31 downto 0);                    -- writedata
			audio_codec_avalon_audio_slave_chipselect       : out std_logic;                                        -- chipselect
			audio_config_avalon_av_config_slave_address     : out std_logic_vector(1 downto 0);                     -- address
			audio_config_avalon_av_config_slave_write       : out std_logic;                                        -- write
			audio_config_avalon_av_config_slave_read        : out std_logic;                                        -- read
			audio_config_avalon_av_config_slave_readdata    : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			audio_config_avalon_av_config_slave_writedata   : out std_logic_vector(31 downto 0);                    -- writedata
			audio_config_avalon_av_config_slave_byteenable  : out std_logic_vector(3 downto 0);                     -- byteenable
			audio_config_avalon_av_config_slave_waitrequest : in  std_logic                     := 'X';             -- waitrequest
			nios2_gen2_0_debug_mem_slave_address            : out std_logic_vector(8 downto 0);                     -- address
			nios2_gen2_0_debug_mem_slave_write              : out std_logic;                                        -- write
			nios2_gen2_0_debug_mem_slave_read               : out std_logic;                                        -- read
			nios2_gen2_0_debug_mem_slave_readdata           : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			nios2_gen2_0_debug_mem_slave_writedata          : out std_logic_vector(31 downto 0);                    -- writedata
			nios2_gen2_0_debug_mem_slave_byteenable         : out std_logic_vector(3 downto 0);                     -- byteenable
			nios2_gen2_0_debug_mem_slave_waitrequest        : in  std_logic                     := 'X';             -- waitrequest
			nios2_gen2_0_debug_mem_slave_debugaccess        : out std_logic;                                        -- debugaccess
			onchip_memory2_0_s1_address                     : out std_logic_vector(16 downto 0);                    -- address
			onchip_memory2_0_s1_write                       : out std_logic;                                        -- write
			onchip_memory2_0_s1_readdata                    : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			onchip_memory2_0_s1_writedata                   : out std_logic_vector(31 downto 0);                    -- writedata
			onchip_memory2_0_s1_byteenable                  : out std_logic_vector(3 downto 0);                     -- byteenable
			onchip_memory2_0_s1_chipselect                  : out std_logic;                                        -- chipselect
			onchip_memory2_0_s1_clken                       : out std_logic;                                        -- clken
			sysid_qsys_0_control_slave_address              : out std_logic_vector(0 downto 0);                     -- address
			sysid_qsys_0_control_slave_readdata             : in  std_logic_vector(31 downto 0) := (others => 'X')  -- readdata
		);
	end component system_mm_interconnect_0;

	component system_irq_mapper is
		port (
			clk           : in  std_logic                     := 'X'; -- clk
			reset         : in  std_logic                     := 'X'; -- reset
			receiver0_irq : in  std_logic                     := 'X'; -- irq
			sender_irq    : out std_logic_vector(31 downto 0)         -- irq
		);
	end component system_irq_mapper;

	component altera_irq_clock_crosser is
		generic (
			IRQ_WIDTH : integer := 1
		);
		port (
			receiver_clk   : in  std_logic                    := 'X';             -- clk
			sender_clk     : in  std_logic                    := 'X';             -- clk
			receiver_reset : in  std_logic                    := 'X';             -- reset
			sender_reset   : in  std_logic                    := 'X';             -- reset
			receiver_irq   : in  std_logic_vector(0 downto 0) := (others => 'X'); -- irq
			sender_irq     : out std_logic_vector(0 downto 0)                     -- irq
		);
	end component altera_irq_clock_crosser;

	component system_rst_controller is
		generic (
			NUM_RESET_INPUTS          : integer := 6;
			OUTPUT_RESET_SYNC_EDGES   : string  := "deassert";
			SYNC_DEPTH                : integer := 2;
			RESET_REQUEST_PRESENT     : integer := 0;
			RESET_REQ_WAIT_TIME       : integer := 1;
			MIN_RST_ASSERTION_TIME    : integer := 3;
			RESET_REQ_EARLY_DSRT_TIME : integer := 1;
			USE_RESET_REQUEST_IN0     : integer := 0;
			USE_RESET_REQUEST_IN1     : integer := 0;
			USE_RESET_REQUEST_IN2     : integer := 0;
			USE_RESET_REQUEST_IN3     : integer := 0;
			USE_RESET_REQUEST_IN4     : integer := 0;
			USE_RESET_REQUEST_IN5     : integer := 0;
			USE_RESET_REQUEST_IN6     : integer := 0;
			USE_RESET_REQUEST_IN7     : integer := 0;
			USE_RESET_REQUEST_IN8     : integer := 0;
			USE_RESET_REQUEST_IN9     : integer := 0;
			USE_RESET_REQUEST_IN10    : integer := 0;
			USE_RESET_REQUEST_IN11    : integer := 0;
			USE_RESET_REQUEST_IN12    : integer := 0;
			USE_RESET_REQUEST_IN13    : integer := 0;
			USE_RESET_REQUEST_IN14    : integer := 0;
			USE_RESET_REQUEST_IN15    : integer := 0;
			ADAPT_RESET_REQUEST       : integer := 0
		);
		port (
			reset_in0      : in  std_logic := 'X'; -- reset_in0.reset
			clk            : in  std_logic := 'X'; --       clk.clk
			reset_out      : out std_logic;        -- reset_out.reset
			reset_in1      : in  std_logic := 'X';
			reset_in10     : in  std_logic := 'X';
			reset_in11     : in  std_logic := 'X';
			reset_in12     : in  std_logic := 'X';
			reset_in13     : in  std_logic := 'X';
			reset_in14     : in  std_logic := 'X';
			reset_in15     : in  std_logic := 'X';
			reset_in2      : in  std_logic := 'X';
			reset_in3      : in  std_logic := 'X';
			reset_in4      : in  std_logic := 'X';
			reset_in5      : in  std_logic := 'X';
			reset_in6      : in  std_logic := 'X';
			reset_in7      : in  std_logic := 'X';
			reset_in8      : in  std_logic := 'X';
			reset_in9      : in  std_logic := 'X';
			reset_req      : out std_logic;
			reset_req_in0  : in  std_logic := 'X';
			reset_req_in1  : in  std_logic := 'X';
			reset_req_in10 : in  std_logic := 'X';
			reset_req_in11 : in  std_logic := 'X';
			reset_req_in12 : in  std_logic := 'X';
			reset_req_in13 : in  std_logic := 'X';
			reset_req_in14 : in  std_logic := 'X';
			reset_req_in15 : in  std_logic := 'X';
			reset_req_in2  : in  std_logic := 'X';
			reset_req_in3  : in  std_logic := 'X';
			reset_req_in4  : in  std_logic := 'X';
			reset_req_in5  : in  std_logic := 'X';
			reset_req_in6  : in  std_logic := 'X';
			reset_req_in7  : in  std_logic := 'X';
			reset_req_in8  : in  std_logic := 'X';
			reset_req_in9  : in  std_logic := 'X'
		);
	end component system_rst_controller;

	component system_rst_controller_001 is
		generic (
			NUM_RESET_INPUTS          : integer := 6;
			OUTPUT_RESET_SYNC_EDGES   : string  := "deassert";
			SYNC_DEPTH                : integer := 2;
			RESET_REQUEST_PRESENT     : integer := 0;
			RESET_REQ_WAIT_TIME       : integer := 1;
			MIN_RST_ASSERTION_TIME    : integer := 3;
			RESET_REQ_EARLY_DSRT_TIME : integer := 1;
			USE_RESET_REQUEST_IN0     : integer := 0;
			USE_RESET_REQUEST_IN1     : integer := 0;
			USE_RESET_REQUEST_IN2     : integer := 0;
			USE_RESET_REQUEST_IN3     : integer := 0;
			USE_RESET_REQUEST_IN4     : integer := 0;
			USE_RESET_REQUEST_IN5     : integer := 0;
			USE_RESET_REQUEST_IN6     : integer := 0;
			USE_RESET_REQUEST_IN7     : integer := 0;
			USE_RESET_REQUEST_IN8     : integer := 0;
			USE_RESET_REQUEST_IN9     : integer := 0;
			USE_RESET_REQUEST_IN10    : integer := 0;
			USE_RESET_REQUEST_IN11    : integer := 0;
			USE_RESET_REQUEST_IN12    : integer := 0;
			USE_RESET_REQUEST_IN13    : integer := 0;
			USE_RESET_REQUEST_IN14    : integer := 0;
			USE_RESET_REQUEST_IN15    : integer := 0;
			ADAPT_RESET_REQUEST       : integer := 0
		);
		port (
			reset_in0      : in  std_logic := 'X'; -- reset_in0.reset
			clk            : in  std_logic := 'X'; --       clk.clk
			reset_out      : out std_logic;        -- reset_out.reset
			reset_req      : out std_logic;        --          .reset_req
			reset_in1      : in  std_logic := 'X';
			reset_in10     : in  std_logic := 'X';
			reset_in11     : in  std_logic := 'X';
			reset_in12     : in  std_logic := 'X';
			reset_in13     : in  std_logic := 'X';
			reset_in14     : in  std_logic := 'X';
			reset_in15     : in  std_logic := 'X';
			reset_in2      : in  std_logic := 'X';
			reset_in3      : in  std_logic := 'X';
			reset_in4      : in  std_logic := 'X';
			reset_in5      : in  std_logic := 'X';
			reset_in6      : in  std_logic := 'X';
			reset_in7      : in  std_logic := 'X';
			reset_in8      : in  std_logic := 'X';
			reset_in9      : in  std_logic := 'X';
			reset_req_in0  : in  std_logic := 'X';
			reset_req_in1  : in  std_logic := 'X';
			reset_req_in10 : in  std_logic := 'X';
			reset_req_in11 : in  std_logic := 'X';
			reset_req_in12 : in  std_logic := 'X';
			reset_req_in13 : in  std_logic := 'X';
			reset_req_in14 : in  std_logic := 'X';
			reset_req_in15 : in  std_logic := 'X';
			reset_req_in2  : in  std_logic := 'X';
			reset_req_in3  : in  std_logic := 'X';
			reset_req_in4  : in  std_logic := 'X';
			reset_req_in5  : in  std_logic := 'X';
			reset_req_in6  : in  std_logic := 'X';
			reset_req_in7  : in  std_logic := 'X';
			reset_req_in8  : in  std_logic := 'X';
			reset_req_in9  : in  std_logic := 'X'
		);
	end component system_rst_controller_001;

	signal audio_pll_0_audio_clk_clk                                         : std_logic;                     -- audio_pll_0:audio_clk_clk -> [audio_pll_1_audio_clk_clk, audio_codec:clk, irq_synchronizer:receiver_clk, mm_interconnect_0:clock_bridge_0_out_clk_clk, rst_controller:clk]
	signal nios2_gen2_0_data_master_readdata                                 : std_logic_vector(31 downto 0); -- mm_interconnect_0:nios2_gen2_0_data_master_readdata -> nios2_gen2_0:d_readdata
	signal nios2_gen2_0_data_master_waitrequest                              : std_logic;                     -- mm_interconnect_0:nios2_gen2_0_data_master_waitrequest -> nios2_gen2_0:d_waitrequest
	signal nios2_gen2_0_data_master_debugaccess                              : std_logic;                     -- nios2_gen2_0:debug_mem_slave_debugaccess_to_roms -> mm_interconnect_0:nios2_gen2_0_data_master_debugaccess
	signal nios2_gen2_0_data_master_address                                  : std_logic_vector(20 downto 0); -- nios2_gen2_0:d_address -> mm_interconnect_0:nios2_gen2_0_data_master_address
	signal nios2_gen2_0_data_master_byteenable                               : std_logic_vector(3 downto 0);  -- nios2_gen2_0:d_byteenable -> mm_interconnect_0:nios2_gen2_0_data_master_byteenable
	signal nios2_gen2_0_data_master_read                                     : std_logic;                     -- nios2_gen2_0:d_read -> mm_interconnect_0:nios2_gen2_0_data_master_read
	signal nios2_gen2_0_data_master_write                                    : std_logic;                     -- nios2_gen2_0:d_write -> mm_interconnect_0:nios2_gen2_0_data_master_write
	signal nios2_gen2_0_data_master_writedata                                : std_logic_vector(31 downto 0); -- nios2_gen2_0:d_writedata -> mm_interconnect_0:nios2_gen2_0_data_master_writedata
	signal nios2_gen2_0_instruction_master_readdata                          : std_logic_vector(31 downto 0); -- mm_interconnect_0:nios2_gen2_0_instruction_master_readdata -> nios2_gen2_0:i_readdata
	signal nios2_gen2_0_instruction_master_waitrequest                       : std_logic;                     -- mm_interconnect_0:nios2_gen2_0_instruction_master_waitrequest -> nios2_gen2_0:i_waitrequest
	signal nios2_gen2_0_instruction_master_address                           : std_logic_vector(20 downto 0); -- nios2_gen2_0:i_address -> mm_interconnect_0:nios2_gen2_0_instruction_master_address
	signal nios2_gen2_0_instruction_master_read                              : std_logic;                     -- nios2_gen2_0:i_read -> mm_interconnect_0:nios2_gen2_0_instruction_master_read
	signal mm_interconnect_0_audio_codec_avalon_audio_slave_chipselect       : std_logic;                     -- mm_interconnect_0:audio_codec_avalon_audio_slave_chipselect -> audio_codec:chipselect
	signal mm_interconnect_0_audio_codec_avalon_audio_slave_readdata         : std_logic_vector(31 downto 0); -- audio_codec:readdata -> mm_interconnect_0:audio_codec_avalon_audio_slave_readdata
	signal mm_interconnect_0_audio_codec_avalon_audio_slave_address          : std_logic_vector(1 downto 0);  -- mm_interconnect_0:audio_codec_avalon_audio_slave_address -> audio_codec:address
	signal mm_interconnect_0_audio_codec_avalon_audio_slave_read             : std_logic;                     -- mm_interconnect_0:audio_codec_avalon_audio_slave_read -> audio_codec:read
	signal mm_interconnect_0_audio_codec_avalon_audio_slave_write            : std_logic;                     -- mm_interconnect_0:audio_codec_avalon_audio_slave_write -> audio_codec:write
	signal mm_interconnect_0_audio_codec_avalon_audio_slave_writedata        : std_logic_vector(31 downto 0); -- mm_interconnect_0:audio_codec_avalon_audio_slave_writedata -> audio_codec:writedata
	signal mm_interconnect_0_audio_config_avalon_av_config_slave_readdata    : std_logic_vector(31 downto 0); -- audio_config:readdata -> mm_interconnect_0:audio_config_avalon_av_config_slave_readdata
	signal mm_interconnect_0_audio_config_avalon_av_config_slave_waitrequest : std_logic;                     -- audio_config:waitrequest -> mm_interconnect_0:audio_config_avalon_av_config_slave_waitrequest
	signal mm_interconnect_0_audio_config_avalon_av_config_slave_address     : std_logic_vector(1 downto 0);  -- mm_interconnect_0:audio_config_avalon_av_config_slave_address -> audio_config:address
	signal mm_interconnect_0_audio_config_avalon_av_config_slave_read        : std_logic;                     -- mm_interconnect_0:audio_config_avalon_av_config_slave_read -> audio_config:read
	signal mm_interconnect_0_audio_config_avalon_av_config_slave_byteenable  : std_logic_vector(3 downto 0);  -- mm_interconnect_0:audio_config_avalon_av_config_slave_byteenable -> audio_config:byteenable
	signal mm_interconnect_0_audio_config_avalon_av_config_slave_write       : std_logic;                     -- mm_interconnect_0:audio_config_avalon_av_config_slave_write -> audio_config:write
	signal mm_interconnect_0_audio_config_avalon_av_config_slave_writedata   : std_logic_vector(31 downto 0); -- mm_interconnect_0:audio_config_avalon_av_config_slave_writedata -> audio_config:writedata
	signal mm_interconnect_0_sysid_qsys_0_control_slave_readdata             : std_logic_vector(31 downto 0); -- sysid_qsys_0:readdata -> mm_interconnect_0:sysid_qsys_0_control_slave_readdata
	signal mm_interconnect_0_sysid_qsys_0_control_slave_address              : std_logic_vector(0 downto 0);  -- mm_interconnect_0:sysid_qsys_0_control_slave_address -> sysid_qsys_0:address
	signal mm_interconnect_0_nios2_gen2_0_debug_mem_slave_readdata           : std_logic_vector(31 downto 0); -- nios2_gen2_0:debug_mem_slave_readdata -> mm_interconnect_0:nios2_gen2_0_debug_mem_slave_readdata
	signal mm_interconnect_0_nios2_gen2_0_debug_mem_slave_waitrequest        : std_logic;                     -- nios2_gen2_0:debug_mem_slave_waitrequest -> mm_interconnect_0:nios2_gen2_0_debug_mem_slave_waitrequest
	signal mm_interconnect_0_nios2_gen2_0_debug_mem_slave_debugaccess        : std_logic;                     -- mm_interconnect_0:nios2_gen2_0_debug_mem_slave_debugaccess -> nios2_gen2_0:debug_mem_slave_debugaccess
	signal mm_interconnect_0_nios2_gen2_0_debug_mem_slave_address            : std_logic_vector(8 downto 0);  -- mm_interconnect_0:nios2_gen2_0_debug_mem_slave_address -> nios2_gen2_0:debug_mem_slave_address
	signal mm_interconnect_0_nios2_gen2_0_debug_mem_slave_read               : std_logic;                     -- mm_interconnect_0:nios2_gen2_0_debug_mem_slave_read -> nios2_gen2_0:debug_mem_slave_read
	signal mm_interconnect_0_nios2_gen2_0_debug_mem_slave_byteenable         : std_logic_vector(3 downto 0);  -- mm_interconnect_0:nios2_gen2_0_debug_mem_slave_byteenable -> nios2_gen2_0:debug_mem_slave_byteenable
	signal mm_interconnect_0_nios2_gen2_0_debug_mem_slave_write              : std_logic;                     -- mm_interconnect_0:nios2_gen2_0_debug_mem_slave_write -> nios2_gen2_0:debug_mem_slave_write
	signal mm_interconnect_0_nios2_gen2_0_debug_mem_slave_writedata          : std_logic_vector(31 downto 0); -- mm_interconnect_0:nios2_gen2_0_debug_mem_slave_writedata -> nios2_gen2_0:debug_mem_slave_writedata
	signal mm_interconnect_0_onchip_memory2_0_s1_chipselect                  : std_logic;                     -- mm_interconnect_0:onchip_memory2_0_s1_chipselect -> onchip_memory2_0:chipselect
	signal mm_interconnect_0_onchip_memory2_0_s1_readdata                    : std_logic_vector(31 downto 0); -- onchip_memory2_0:readdata -> mm_interconnect_0:onchip_memory2_0_s1_readdata
	signal mm_interconnect_0_onchip_memory2_0_s1_address                     : std_logic_vector(16 downto 0); -- mm_interconnect_0:onchip_memory2_0_s1_address -> onchip_memory2_0:address
	signal mm_interconnect_0_onchip_memory2_0_s1_byteenable                  : std_logic_vector(3 downto 0);  -- mm_interconnect_0:onchip_memory2_0_s1_byteenable -> onchip_memory2_0:byteenable
	signal mm_interconnect_0_onchip_memory2_0_s1_write                       : std_logic;                     -- mm_interconnect_0:onchip_memory2_0_s1_write -> onchip_memory2_0:write
	signal mm_interconnect_0_onchip_memory2_0_s1_writedata                   : std_logic_vector(31 downto 0); -- mm_interconnect_0:onchip_memory2_0_s1_writedata -> onchip_memory2_0:writedata
	signal mm_interconnect_0_onchip_memory2_0_s1_clken                       : std_logic;                     -- mm_interconnect_0:onchip_memory2_0_s1_clken -> onchip_memory2_0:clken
	signal nios2_gen2_0_irq_irq                                              : std_logic_vector(31 downto 0); -- irq_mapper:sender_irq -> nios2_gen2_0:irq
	signal irq_mapper_receiver0_irq                                          : std_logic;                     -- irq_synchronizer:sender_irq -> irq_mapper:receiver0_irq
	signal irq_synchronizer_receiver_irq                                     : std_logic_vector(0 downto 0);  -- audio_codec:irq -> irq_synchronizer:receiver_irq
	signal rst_controller_reset_out_reset                                    : std_logic;                     -- rst_controller:reset_out -> [audio_codec:reset, irq_synchronizer:receiver_reset, mm_interconnect_0:audio_codec_reset_reset_bridge_in_reset_reset]
	signal rst_controller_001_reset_out_reset                                : std_logic;                     -- rst_controller_001:reset_out -> [audio_config:reset, irq_mapper:reset, irq_synchronizer:sender_reset, mm_interconnect_0:nios2_gen2_0_reset_reset_bridge_in_reset_reset, onchip_memory2_0:reset, rst_controller_001_reset_out_reset:in, rst_translator:in_reset]
	signal rst_controller_001_reset_out_reset_req                            : std_logic;                     -- rst_controller_001:reset_req -> [nios2_gen2_0:reset_req, onchip_memory2_0:reset_req, rst_translator:reset_req_in]
	signal reset_reset_n_ports_inv                                           : std_logic;                     -- reset_reset_n:inv -> [audio_pll_0:ref_reset_reset, rst_controller:reset_in0, rst_controller_001:reset_in0]
	signal rst_controller_001_reset_out_reset_ports_inv                      : std_logic;                     -- rst_controller_001_reset_out_reset:inv -> [nios2_gen2_0:reset_n, sysid_qsys_0:reset_n]

begin

	audio_codec : component system_audio_codec
		port map (
			clk         => audio_pll_0_audio_clk_clk,                                   --                clk.clk
			reset       => rst_controller_reset_out_reset,                              --              reset.reset
			address     => mm_interconnect_0_audio_codec_avalon_audio_slave_address,    -- avalon_audio_slave.address
			chipselect  => mm_interconnect_0_audio_codec_avalon_audio_slave_chipselect, --                   .chipselect
			read        => mm_interconnect_0_audio_codec_avalon_audio_slave_read,       --                   .read
			write       => mm_interconnect_0_audio_codec_avalon_audio_slave_write,      --                   .write
			writedata   => mm_interconnect_0_audio_codec_avalon_audio_slave_writedata,  --                   .writedata
			readdata    => mm_interconnect_0_audio_codec_avalon_audio_slave_readdata,   --                   .readdata
			irq         => irq_synchronizer_receiver_irq(0),                            --          interrupt.irq
			AUD_ADCDAT  => audio_codec_external_interface_ADCDAT,                       -- external_interface.export
			AUD_ADCLRCK => audio_codec_external_interface_ADCLRCK,                      --                   .export
			AUD_BCLK    => audio_codec_external_interface_BCLK,                         --                   .export
			AUD_DACDAT  => audio_codec_external_interface_DACDAT,                       --                   .export
			AUD_DACLRCK => audio_codec_external_interface_DACLRCK                       --                   .export
		);

	audio_config : component system_audio_config
		port map (
			clk         => clk_clk,                                                           --                    clk.clk
			reset       => rst_controller_001_reset_out_reset,                                --                  reset.reset
			address     => mm_interconnect_0_audio_config_avalon_av_config_slave_address,     -- avalon_av_config_slave.address
			byteenable  => mm_interconnect_0_audio_config_avalon_av_config_slave_byteenable,  --                       .byteenable
			read        => mm_interconnect_0_audio_config_avalon_av_config_slave_read,        --                       .read
			write       => mm_interconnect_0_audio_config_avalon_av_config_slave_write,       --                       .write
			writedata   => mm_interconnect_0_audio_config_avalon_av_config_slave_writedata,   --                       .writedata
			readdata    => mm_interconnect_0_audio_config_avalon_av_config_slave_readdata,    --                       .readdata
			waitrequest => mm_interconnect_0_audio_config_avalon_av_config_slave_waitrequest, --                       .waitrequest
			I2C_SDAT    => audio_config_external_interface_SDAT,                              --     external_interface.export
			I2C_SCLK    => audio_config_external_interface_SCLK                               --                       .export
		);

	audio_pll_0 : component system_audio_pll_0
		port map (
			ref_clk_clk        => clk_clk,                   --      ref_clk.clk
			ref_reset_reset    => reset_reset_n_ports_inv,   --    ref_reset.reset
			audio_clk_clk      => audio_pll_0_audio_clk_clk, --    audio_clk.clk
			reset_source_reset => open                       -- reset_source.reset
		);

	nios2_gen2_0 : component system_nios2_gen2_0
		port map (
			clk                                 => clk_clk,                                                    --                       clk.clk
			reset_n                             => rst_controller_001_reset_out_reset_ports_inv,               --                     reset.reset_n
			reset_req                           => rst_controller_001_reset_out_reset_req,                     --                          .reset_req
			d_address                           => nios2_gen2_0_data_master_address,                           --               data_master.address
			d_byteenable                        => nios2_gen2_0_data_master_byteenable,                        --                          .byteenable
			d_read                              => nios2_gen2_0_data_master_read,                              --                          .read
			d_readdata                          => nios2_gen2_0_data_master_readdata,                          --                          .readdata
			d_waitrequest                       => nios2_gen2_0_data_master_waitrequest,                       --                          .waitrequest
			d_write                             => nios2_gen2_0_data_master_write,                             --                          .write
			d_writedata                         => nios2_gen2_0_data_master_writedata,                         --                          .writedata
			debug_mem_slave_debugaccess_to_roms => nios2_gen2_0_data_master_debugaccess,                       --                          .debugaccess
			i_address                           => nios2_gen2_0_instruction_master_address,                    --        instruction_master.address
			i_read                              => nios2_gen2_0_instruction_master_read,                       --                          .read
			i_readdata                          => nios2_gen2_0_instruction_master_readdata,                   --                          .readdata
			i_waitrequest                       => nios2_gen2_0_instruction_master_waitrequest,                --                          .waitrequest
			irq                                 => nios2_gen2_0_irq_irq,                                       --                       irq.irq
			debug_reset_request                 => open,                                                       --       debug_reset_request.reset
			debug_mem_slave_address             => mm_interconnect_0_nios2_gen2_0_debug_mem_slave_address,     --           debug_mem_slave.address
			debug_mem_slave_byteenable          => mm_interconnect_0_nios2_gen2_0_debug_mem_slave_byteenable,  --                          .byteenable
			debug_mem_slave_debugaccess         => mm_interconnect_0_nios2_gen2_0_debug_mem_slave_debugaccess, --                          .debugaccess
			debug_mem_slave_read                => mm_interconnect_0_nios2_gen2_0_debug_mem_slave_read,        --                          .read
			debug_mem_slave_readdata            => mm_interconnect_0_nios2_gen2_0_debug_mem_slave_readdata,    --                          .readdata
			debug_mem_slave_waitrequest         => mm_interconnect_0_nios2_gen2_0_debug_mem_slave_waitrequest, --                          .waitrequest
			debug_mem_slave_write               => mm_interconnect_0_nios2_gen2_0_debug_mem_slave_write,       --                          .write
			debug_mem_slave_writedata           => mm_interconnect_0_nios2_gen2_0_debug_mem_slave_writedata,   --                          .writedata
			dummy_ci_port                       => open                                                        -- custom_instruction_master.readra
		);

	onchip_memory2_0 : component system_onchip_memory2_0
		port map (
			clk        => clk_clk,                                          --   clk1.clk
			address    => mm_interconnect_0_onchip_memory2_0_s1_address,    --     s1.address
			clken      => mm_interconnect_0_onchip_memory2_0_s1_clken,      --       .clken
			chipselect => mm_interconnect_0_onchip_memory2_0_s1_chipselect, --       .chipselect
			write      => mm_interconnect_0_onchip_memory2_0_s1_write,      --       .write
			readdata   => mm_interconnect_0_onchip_memory2_0_s1_readdata,   --       .readdata
			writedata  => mm_interconnect_0_onchip_memory2_0_s1_writedata,  --       .writedata
			byteenable => mm_interconnect_0_onchip_memory2_0_s1_byteenable, --       .byteenable
			reset      => rst_controller_001_reset_out_reset,               -- reset1.reset
			reset_req  => rst_controller_001_reset_out_reset_req,           --       .reset_req
			freeze     => '0'                                               -- (terminated)
		);

	sysid_qsys_0 : component system_sysid_qsys_0
		port map (
			clock    => clk_clk,                                                 --           clk.clk
			reset_n  => rst_controller_001_reset_out_reset_ports_inv,            --         reset.reset_n
			readdata => mm_interconnect_0_sysid_qsys_0_control_slave_readdata,   -- control_slave.readdata
			address  => mm_interconnect_0_sysid_qsys_0_control_slave_address(0)  --              .address
		);

	mm_interconnect_0 : component system_mm_interconnect_0
		port map (
			clk_0_clk_clk                                   => clk_clk,                                                           --                                clk_0_clk.clk
			clock_bridge_0_out_clk_clk                      => audio_pll_0_audio_clk_clk,                                         --                   clock_bridge_0_out_clk.clk
			audio_codec_reset_reset_bridge_in_reset_reset   => rst_controller_reset_out_reset,                                    --  audio_codec_reset_reset_bridge_in_reset.reset
			nios2_gen2_0_reset_reset_bridge_in_reset_reset  => rst_controller_001_reset_out_reset,                                -- nios2_gen2_0_reset_reset_bridge_in_reset.reset
			nios2_gen2_0_data_master_address                => nios2_gen2_0_data_master_address,                                  --                 nios2_gen2_0_data_master.address
			nios2_gen2_0_data_master_waitrequest            => nios2_gen2_0_data_master_waitrequest,                              --                                         .waitrequest
			nios2_gen2_0_data_master_byteenable             => nios2_gen2_0_data_master_byteenable,                               --                                         .byteenable
			nios2_gen2_0_data_master_read                   => nios2_gen2_0_data_master_read,                                     --                                         .read
			nios2_gen2_0_data_master_readdata               => nios2_gen2_0_data_master_readdata,                                 --                                         .readdata
			nios2_gen2_0_data_master_write                  => nios2_gen2_0_data_master_write,                                    --                                         .write
			nios2_gen2_0_data_master_writedata              => nios2_gen2_0_data_master_writedata,                                --                                         .writedata
			nios2_gen2_0_data_master_debugaccess            => nios2_gen2_0_data_master_debugaccess,                              --                                         .debugaccess
			nios2_gen2_0_instruction_master_address         => nios2_gen2_0_instruction_master_address,                           --          nios2_gen2_0_instruction_master.address
			nios2_gen2_0_instruction_master_waitrequest     => nios2_gen2_0_instruction_master_waitrequest,                       --                                         .waitrequest
			nios2_gen2_0_instruction_master_read            => nios2_gen2_0_instruction_master_read,                              --                                         .read
			nios2_gen2_0_instruction_master_readdata        => nios2_gen2_0_instruction_master_readdata,                          --                                         .readdata
			audio_codec_avalon_audio_slave_address          => mm_interconnect_0_audio_codec_avalon_audio_slave_address,          --           audio_codec_avalon_audio_slave.address
			audio_codec_avalon_audio_slave_write            => mm_interconnect_0_audio_codec_avalon_audio_slave_write,            --                                         .write
			audio_codec_avalon_audio_slave_read             => mm_interconnect_0_audio_codec_avalon_audio_slave_read,             --                                         .read
			audio_codec_avalon_audio_slave_readdata         => mm_interconnect_0_audio_codec_avalon_audio_slave_readdata,         --                                         .readdata
			audio_codec_avalon_audio_slave_writedata        => mm_interconnect_0_audio_codec_avalon_audio_slave_writedata,        --                                         .writedata
			audio_codec_avalon_audio_slave_chipselect       => mm_interconnect_0_audio_codec_avalon_audio_slave_chipselect,       --                                         .chipselect
			audio_config_avalon_av_config_slave_address     => mm_interconnect_0_audio_config_avalon_av_config_slave_address,     --      audio_config_avalon_av_config_slave.address
			audio_config_avalon_av_config_slave_write       => mm_interconnect_0_audio_config_avalon_av_config_slave_write,       --                                         .write
			audio_config_avalon_av_config_slave_read        => mm_interconnect_0_audio_config_avalon_av_config_slave_read,        --                                         .read
			audio_config_avalon_av_config_slave_readdata    => mm_interconnect_0_audio_config_avalon_av_config_slave_readdata,    --                                         .readdata
			audio_config_avalon_av_config_slave_writedata   => mm_interconnect_0_audio_config_avalon_av_config_slave_writedata,   --                                         .writedata
			audio_config_avalon_av_config_slave_byteenable  => mm_interconnect_0_audio_config_avalon_av_config_slave_byteenable,  --                                         .byteenable
			audio_config_avalon_av_config_slave_waitrequest => mm_interconnect_0_audio_config_avalon_av_config_slave_waitrequest, --                                         .waitrequest
			nios2_gen2_0_debug_mem_slave_address            => mm_interconnect_0_nios2_gen2_0_debug_mem_slave_address,            --             nios2_gen2_0_debug_mem_slave.address
			nios2_gen2_0_debug_mem_slave_write              => mm_interconnect_0_nios2_gen2_0_debug_mem_slave_write,              --                                         .write
			nios2_gen2_0_debug_mem_slave_read               => mm_interconnect_0_nios2_gen2_0_debug_mem_slave_read,               --                                         .read
			nios2_gen2_0_debug_mem_slave_readdata           => mm_interconnect_0_nios2_gen2_0_debug_mem_slave_readdata,           --                                         .readdata
			nios2_gen2_0_debug_mem_slave_writedata          => mm_interconnect_0_nios2_gen2_0_debug_mem_slave_writedata,          --                                         .writedata
			nios2_gen2_0_debug_mem_slave_byteenable         => mm_interconnect_0_nios2_gen2_0_debug_mem_slave_byteenable,         --                                         .byteenable
			nios2_gen2_0_debug_mem_slave_waitrequest        => mm_interconnect_0_nios2_gen2_0_debug_mem_slave_waitrequest,        --                                         .waitrequest
			nios2_gen2_0_debug_mem_slave_debugaccess        => mm_interconnect_0_nios2_gen2_0_debug_mem_slave_debugaccess,        --                                         .debugaccess
			onchip_memory2_0_s1_address                     => mm_interconnect_0_onchip_memory2_0_s1_address,                     --                      onchip_memory2_0_s1.address
			onchip_memory2_0_s1_write                       => mm_interconnect_0_onchip_memory2_0_s1_write,                       --                                         .write
			onchip_memory2_0_s1_readdata                    => mm_interconnect_0_onchip_memory2_0_s1_readdata,                    --                                         .readdata
			onchip_memory2_0_s1_writedata                   => mm_interconnect_0_onchip_memory2_0_s1_writedata,                   --                                         .writedata
			onchip_memory2_0_s1_byteenable                  => mm_interconnect_0_onchip_memory2_0_s1_byteenable,                  --                                         .byteenable
			onchip_memory2_0_s1_chipselect                  => mm_interconnect_0_onchip_memory2_0_s1_chipselect,                  --                                         .chipselect
			onchip_memory2_0_s1_clken                       => mm_interconnect_0_onchip_memory2_0_s1_clken,                       --                                         .clken
			sysid_qsys_0_control_slave_address              => mm_interconnect_0_sysid_qsys_0_control_slave_address,              --               sysid_qsys_0_control_slave.address
			sysid_qsys_0_control_slave_readdata             => mm_interconnect_0_sysid_qsys_0_control_slave_readdata              --                                         .readdata
		);

	irq_mapper : component system_irq_mapper
		port map (
			clk           => clk_clk,                            --       clk.clk
			reset         => rst_controller_001_reset_out_reset, -- clk_reset.reset
			receiver0_irq => irq_mapper_receiver0_irq,           -- receiver0.irq
			sender_irq    => nios2_gen2_0_irq_irq                --    sender.irq
		);

	irq_synchronizer : component altera_irq_clock_crosser
		generic map (
			IRQ_WIDTH => 1
		)
		port map (
			receiver_clk   => audio_pll_0_audio_clk_clk,          --       receiver_clk.clk
			sender_clk     => clk_clk,                            --         sender_clk.clk
			receiver_reset => rst_controller_reset_out_reset,     -- receiver_clk_reset.reset
			sender_reset   => rst_controller_001_reset_out_reset, --   sender_clk_reset.reset
			receiver_irq   => irq_synchronizer_receiver_irq,      --           receiver.irq
			sender_irq(0)  => irq_mapper_receiver0_irq            --             sender.irq
		);

	rst_controller : component system_rst_controller
		generic map (
			NUM_RESET_INPUTS          => 1,
			OUTPUT_RESET_SYNC_EDGES   => "deassert",
			SYNC_DEPTH                => 2,
			RESET_REQUEST_PRESENT     => 0,
			RESET_REQ_WAIT_TIME       => 1,
			MIN_RST_ASSERTION_TIME    => 3,
			RESET_REQ_EARLY_DSRT_TIME => 1,
			USE_RESET_REQUEST_IN0     => 0,
			USE_RESET_REQUEST_IN1     => 0,
			USE_RESET_REQUEST_IN2     => 0,
			USE_RESET_REQUEST_IN3     => 0,
			USE_RESET_REQUEST_IN4     => 0,
			USE_RESET_REQUEST_IN5     => 0,
			USE_RESET_REQUEST_IN6     => 0,
			USE_RESET_REQUEST_IN7     => 0,
			USE_RESET_REQUEST_IN8     => 0,
			USE_RESET_REQUEST_IN9     => 0,
			USE_RESET_REQUEST_IN10    => 0,
			USE_RESET_REQUEST_IN11    => 0,
			USE_RESET_REQUEST_IN12    => 0,
			USE_RESET_REQUEST_IN13    => 0,
			USE_RESET_REQUEST_IN14    => 0,
			USE_RESET_REQUEST_IN15    => 0,
			ADAPT_RESET_REQUEST       => 0
		)
		port map (
			reset_in0      => reset_reset_n_ports_inv,        -- reset_in0.reset
			clk            => audio_pll_0_audio_clk_clk,      --       clk.clk
			reset_out      => rst_controller_reset_out_reset, -- reset_out.reset
			reset_req      => open,                           -- (terminated)
			reset_req_in0  => '0',                            -- (terminated)
			reset_in1      => '0',                            -- (terminated)
			reset_req_in1  => '0',                            -- (terminated)
			reset_in2      => '0',                            -- (terminated)
			reset_req_in2  => '0',                            -- (terminated)
			reset_in3      => '0',                            -- (terminated)
			reset_req_in3  => '0',                            -- (terminated)
			reset_in4      => '0',                            -- (terminated)
			reset_req_in4  => '0',                            -- (terminated)
			reset_in5      => '0',                            -- (terminated)
			reset_req_in5  => '0',                            -- (terminated)
			reset_in6      => '0',                            -- (terminated)
			reset_req_in6  => '0',                            -- (terminated)
			reset_in7      => '0',                            -- (terminated)
			reset_req_in7  => '0',                            -- (terminated)
			reset_in8      => '0',                            -- (terminated)
			reset_req_in8  => '0',                            -- (terminated)
			reset_in9      => '0',                            -- (terminated)
			reset_req_in9  => '0',                            -- (terminated)
			reset_in10     => '0',                            -- (terminated)
			reset_req_in10 => '0',                            -- (terminated)
			reset_in11     => '0',                            -- (terminated)
			reset_req_in11 => '0',                            -- (terminated)
			reset_in12     => '0',                            -- (terminated)
			reset_req_in12 => '0',                            -- (terminated)
			reset_in13     => '0',                            -- (terminated)
			reset_req_in13 => '0',                            -- (terminated)
			reset_in14     => '0',                            -- (terminated)
			reset_req_in14 => '0',                            -- (terminated)
			reset_in15     => '0',                            -- (terminated)
			reset_req_in15 => '0'                             -- (terminated)
		);

	rst_controller_001 : component system_rst_controller_001
		generic map (
			NUM_RESET_INPUTS          => 1,
			OUTPUT_RESET_SYNC_EDGES   => "deassert",
			SYNC_DEPTH                => 2,
			RESET_REQUEST_PRESENT     => 1,
			RESET_REQ_WAIT_TIME       => 1,
			MIN_RST_ASSERTION_TIME    => 3,
			RESET_REQ_EARLY_DSRT_TIME => 1,
			USE_RESET_REQUEST_IN0     => 0,
			USE_RESET_REQUEST_IN1     => 0,
			USE_RESET_REQUEST_IN2     => 0,
			USE_RESET_REQUEST_IN3     => 0,
			USE_RESET_REQUEST_IN4     => 0,
			USE_RESET_REQUEST_IN5     => 0,
			USE_RESET_REQUEST_IN6     => 0,
			USE_RESET_REQUEST_IN7     => 0,
			USE_RESET_REQUEST_IN8     => 0,
			USE_RESET_REQUEST_IN9     => 0,
			USE_RESET_REQUEST_IN10    => 0,
			USE_RESET_REQUEST_IN11    => 0,
			USE_RESET_REQUEST_IN12    => 0,
			USE_RESET_REQUEST_IN13    => 0,
			USE_RESET_REQUEST_IN14    => 0,
			USE_RESET_REQUEST_IN15    => 0,
			ADAPT_RESET_REQUEST       => 0
		)
		port map (
			reset_in0      => reset_reset_n_ports_inv,                -- reset_in0.reset
			clk            => clk_clk,                                --       clk.clk
			reset_out      => rst_controller_001_reset_out_reset,     -- reset_out.reset
			reset_req      => rst_controller_001_reset_out_reset_req, --          .reset_req
			reset_req_in0  => '0',                                    -- (terminated)
			reset_in1      => '0',                                    -- (terminated)
			reset_req_in1  => '0',                                    -- (terminated)
			reset_in2      => '0',                                    -- (terminated)
			reset_req_in2  => '0',                                    -- (terminated)
			reset_in3      => '0',                                    -- (terminated)
			reset_req_in3  => '0',                                    -- (terminated)
			reset_in4      => '0',                                    -- (terminated)
			reset_req_in4  => '0',                                    -- (terminated)
			reset_in5      => '0',                                    -- (terminated)
			reset_req_in5  => '0',                                    -- (terminated)
			reset_in6      => '0',                                    -- (terminated)
			reset_req_in6  => '0',                                    -- (terminated)
			reset_in7      => '0',                                    -- (terminated)
			reset_req_in7  => '0',                                    -- (terminated)
			reset_in8      => '0',                                    -- (terminated)
			reset_req_in8  => '0',                                    -- (terminated)
			reset_in9      => '0',                                    -- (terminated)
			reset_req_in9  => '0',                                    -- (terminated)
			reset_in10     => '0',                                    -- (terminated)
			reset_req_in10 => '0',                                    -- (terminated)
			reset_in11     => '0',                                    -- (terminated)
			reset_req_in11 => '0',                                    -- (terminated)
			reset_in12     => '0',                                    -- (terminated)
			reset_req_in12 => '0',                                    -- (terminated)
			reset_in13     => '0',                                    -- (terminated)
			reset_req_in13 => '0',                                    -- (terminated)
			reset_in14     => '0',                                    -- (terminated)
			reset_req_in14 => '0',                                    -- (terminated)
			reset_in15     => '0',                                    -- (terminated)
			reset_req_in15 => '0'                                     -- (terminated)
		);

	reset_reset_n_ports_inv <= not reset_reset_n;

	rst_controller_001_reset_out_reset_ports_inv <= not rst_controller_001_reset_out_reset;

	audio_pll_1_audio_clk_clk <= audio_pll_0_audio_clk_clk;

end architecture rtl; -- of system
